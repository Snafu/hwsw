yCbCrMUL_inst : yCbCrMUL PORT MAP (
		clock0	 => clock0_sig,
		dataa_0	 => dataa_0_sig,
		dataa_1	 => dataa_1_sig,
		dataa_2	 => dataa_2_sig,
		datab_0	 => datab_0_sig,
		datab_1	 => datab_1_sig,
		datab_2	 => datab_2_sig,
		result	 => result_sig
	);
